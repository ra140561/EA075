LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MAIN IS
PORT(	IN_KEYBOARD:	IN STD_LOGIC_VECTOR(16 DOWNTO 0);
	OUT_ASCII:	BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0);
	OUT_CRIP, OUT_DESC:	BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0));
END MAIN;

ARCHITECTURE Parte4_Behavior OF MAIN IS

	COMPONENT Somador8b IS
	PORT (	a, b:	in std_logic_vector(7 DOWNTO 0);
		cin: 	in std_logic;
		s:	out std_logic_vector(7 downto 0);
		cout: 	out std_logic);
	END COMPONENT;

	COMPONENT Decode IS
	PORT (	IN_KEYBOARD:	in std_logic_vector(16 downto 0);
		OUT_KEY:	out std_logic_vector(7 downto 0));
	END COMPONENT;

	COMPONENT CRIPT IS
	PORT (	IN_CHAR, CRIPT_CHAR:	in std_logic_vector(7 downto 0);
		ENABLE:			in std_logic;
		OUT_CHAR:		out std_logic_vector(7 downto 0));
	END COMPONENT;

	SIGNAL A: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL SPACE: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL IS_SPACE: STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
	SIGNAL OUT_KEY0, OUT_KEY1: STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL FIM: STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '1');

	SIGNAL COUNT: INTEGER RANGE -1 TO 4 := -1;
	SIGNAL CRIPT_CHAR: STD_LOGIC_VECTOR(7 DOWNTO 0) := "01000011";

	SIGNAL 	C_OUT0, C_OUT1: STD_LOGIC := '0';

	SIGNAL ENABLE_C: STD_LOGIC := '1';

BEGIN

	A <= "01000001"; --registrador do valor do caractere 'A' em ASCII
	SPACE <= "00100000"; --registrador do valor do caractere ' ' (space) em ASCII

	DEC: DECODE PORT MAP(IN_KEYBOARD, OUT_KEY0);

	ADD_Q: SOMADOR8B PORT MAP(OUT_KEY0, A, '0', OUT_KEY1, C_OUT1);

	IS_SPACE <= (OTHERS => ((NOT IN_KEYBOARD(16)) AND IN_KEYBOARD(10)));
	
	PROCESS (IN_KEYBOARD)
	BEGIN
		--SELECIONA A CHAVE CRIPTOGRAFADORA
		CASE (COUNT) IS
			WHEN -1 => CRIPT_CHAR <= "01000011"; --C
			WHEN 0 => CRIPT_CHAR <= "01000011"; --C
			WHEN 1 => CRIPT_CHAR <= "01001111"; --O
			WHEN 2 => CRIPT_CHAR <= "01001100"; --L
			WHEN 3 => CRIPT_CHAR <= "01001111"; --O
			WHEN 4 => CRIPT_CHAR <= "01010010"; --R 
			
		END CASE;

		IF((IN_KEYBOARD(16) AND IN_KEYBOARD(15)) = '1') THEN --SE A TECLA "FIM" FOI PRESSIONADA
			FIM <= (OTHERS => '0');				--NADA SERA IMPRESSO
			ENABLE_C <= '0';
		END IF;

		IF(COUNT = 4) THEN 
			COUNT <= 0;
		ELSE
			COUNT <= COUNT + 1;
		END IF;

		IF((IN_KEYBOARD(16) AND IN_KEYBOARD(14)) = '1') THEN--A TECLA 14 SERA A A TECLA RESET
			FIM <= (OTHERS => '1');	
			COUNT <= 0;
			ENABLE_C <= '1';
		END IF;

	END PROCESS;

	OUT_ASCII <= (((NOT IS_SPACE) AND OUT_KEY1) OR (IS_SPACE AND SPACE)) AND FIM;--CONDICOES PARA IMPRESSAO
	CRIPTOGRAFADOR:		CRIPT PORT MAP (OUT_ASCII, CRIPT_CHAR, ENABLE_C, OUT_CRIP);
	DESCRIPTOGRAFADOR:	CRIPT PORT MAP (OUT_CRIP, CRIPT_CHAR, ENABLE_C, OUT_DESC); 

end Parte4_Behavior;
