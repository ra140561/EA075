LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Parte2 IS
PORT(	IN_KEYBOARD:	IN STD_LOGIC_VECTOR(16 DOWNTO 0);
	OUT_ASCII:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END Parte2;

ARCHITECTURE Parte2_Behavior OF Parte2 IS

	COMPONENT Somador8b IS
	PORT (	a, b:	in std_logic_vector(7 DOWNTO 0);
		cin: 	in std_logic;
		s:	out std_logic_vector(7 downto 0);
		cout: 	out std_logic);
	END COMPONENT;

	SIGNAL A: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL Q_A: STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL SPACE: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL OUT_KEY: STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
	SIGNAL OUT_KEY0, OUT_KEY1: STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL IN_BEF: STD_LOGIC_VECTOR(16 DOWNTO 0) := (OTHERS => '0');

	SIGNAL 	C_OUT0, C_OUT1: STD_LOGIC := '0';

	SIGNAL OP: STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL SOM: STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');


BEGIN

	A <= "01000001"; --registrador do valor do caractere 'A' em ASCII
	SPACE <= "00100000"; --registrador do valor do caractere ' ' (space) em ASCII
	
	

	PROCESS (IN_KEYBOARD)
	BEGIN
		
		OP(0) <= NOT IN_KEYBOARD(0);
		OP(1) <= (NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1));
		OP(2) <= ((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2));
		OP(3) <= (((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3));
		OP(4) <= ((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4));
		OP(5) <= (((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5));
		OP(6) <= ((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6));
		OP(7) <= (((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7));
		OP(8) <= ((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8));
		OP(9) <= (((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9));
		OP(10) <= ((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
			 AND (NOT IN_KEYBOARD(10));
		OP(11) <= (((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
			 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11));
		OP(12) <= ((((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
			 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11))) AND (NOT IN_KEYBOARD(12));
		OP(13) <= (((((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
			 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11))) AND (NOT IN_KEYBOARD(12))) AND (NOT IN_KEYBOARD(13));
		OP(14) <= ((((((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
			 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11))) AND (NOT IN_KEYBOARD(12))) AND (NOT IN_KEYBOARD(13))) AND (NOT IN_KEYBOARD(14));
		OP(15) <= (((((((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
			 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
			 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11))) AND (NOT IN_KEYBOARD(12))) AND (NOT IN_KEYBOARD(13))) AND (NOT IN_KEYBOARD(14)))
			 AND (NOT IN_KEYBOARD(15));



		SOM(0) <= (((OP(0) XOR OP(1)) XOR (OP(2) XOR OP(3))) XOR ((OP(4) XOR OP(5)) XOR (OP(6) XOR OP(7))))
			XOR (((OP(8) XOR OP(9)) XOR (OP(10) XOR OP(11))) XOR ((OP(12) XOR OP(13)) XOR (OP(14) XOR OP(15))));
		SOM(1) <= (OP(1) XOR OP(3)) OR (OP(5) XOR OP(7)) OR (OP(9) XOR OP(11)) OR (OP(13) XOR OP(15));
			SOM(2) <= (OP(3) XOR OP(7)) OR (OP(11) XOR OP(15));
		SOM(3) <= OP(7) XOR OP(15);
		SOM(4) <= OP(15);

		IF(IN_BEF(16) = '1') THEN --OUT_KEY RECEBE O RESULTADO DA SOMA DO VALOR DE "A" COM A VARIAVEL SOM
			OUT_KEY <= OUT_KEY0;
		ELSIF(((NOT IN_BEF(16)) AND (NOT IN_BEF(15))) = '1') THEN --SE O BOTAO NAO ESTIVER PRESSIONADO 
			OUT_KEY <= OUT_KEY1;				--E O BOTAO "FIM" TAMBEM N�O 
		END IF;

		IF(((NOT IN_BEF(16)) AND IN_BEF(10)) = '1') THEN --SE A TECLA SPC FOR PRESSIONADA 
			OUT_KEY <= SPACE;					--O REGISTRADOR RECEBE O VALOR DE SPACE
		END IF;

		IF(((NOT IN_KEYBOARD(16)) AND IN_KEYBOARD(15)) = '1') THEN --SE A TECLA "FIM" FOI PRESSIONADA DEVE-SE IMPRIMIR
			OUT_ASCII <= OUT_KEY;					--NA TELA A LETRA ARMAZENADO
		ELSE
			IN_BEF <= IN_KEYBOARD;
		END IF;
	
		

	END PROCESS;
	
	Q_A(4) <= NOT IN_KEYBOARD(16);
	
	ADD_SOM: SOMADOR8B PORT MAP("01000001", SOM, '0', OUT_KEY0, C_OUT0);

	ADD_Q: SOMADOR8B PORT MAP(OUT_KEY0, Q_A, '0', OUT_KEY1, C_OUT1);

end Parte2_Behavior;
