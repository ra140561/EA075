LIBRARY ieee;
USE ieee.std_logic_1164.all;

-- Decodificador do teclado.

ENTITY DECODE IS
PORT (	IN_KEYBOARD:	in std_logic_vector(16 downto 0);
	OUT_KEY:	out std_logic_vector(7 downto 0));
END DECODE;

ARCHITECTURE DECODING OF DECODE IS

COMPONENT Somador8b IS
	PORT (	a, b:	in std_logic_vector(7 DOWNTO 0);
		cin: 	in std_logic;
		s:	out std_logic_vector(7 downto 0);
		cout: 	out std_logic);
	END COMPONENT;

SIGNAL OP: STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
SIGNAL Q_A, SOM: STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
SIGNAL C_OUT: STD_LOGIC;

BEGIN

	OP(0) <= NOT IN_KEYBOARD(0);
	OP(1) <= (NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1));
	OP(2) <= ((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2));
	OP(3) <= (((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3));
	OP(4) <= ((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4));
	OP(5) <= (((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5));
	OP(6) <= ((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6));
	OP(7) <= (((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7));
	OP(8) <= ((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8));
	OP(9) <= (((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9));
	OP(10) <= ((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
		 AND (NOT IN_KEYBOARD(10));
	OP(11) <= (((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
		 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11));
	OP(12) <= ((((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
		 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11))) AND (NOT IN_KEYBOARD(12));
	OP(13) <= (((((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
		 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11))) AND (NOT IN_KEYBOARD(12))) AND (NOT IN_KEYBOARD(13));
	OP(14) <= ((((((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
		 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11))) AND (NOT IN_KEYBOARD(12))) AND (NOT IN_KEYBOARD(13))) AND (NOT IN_KEYBOARD(14));
	OP(15) <= (((((((((((((((NOT IN_KEYBOARD(0)) AND (NOT IN_KEYBOARD(1))) AND (NOT IN_KEYBOARD(2))) AND (NOT IN_KEYBOARD(3))) AND (NOT IN_KEYBOARD(4)))
		 AND (NOT IN_KEYBOARD(5))) AND (NOT IN_KEYBOARD(6))) AND (NOT IN_KEYBOARD(7))) AND (NOT IN_KEYBOARD(8))) AND (NOT IN_KEYBOARD(9)))
		 AND (NOT IN_KEYBOARD(10))) AND (NOT IN_KEYBOARD(11))) AND (NOT IN_KEYBOARD(12))) AND (NOT IN_KEYBOARD(13))) AND (NOT IN_KEYBOARD(14)))
		 AND (NOT IN_KEYBOARD(15));

	SOM(0) <= (((OP(0) XOR OP(1)) XOR (OP(2) XOR OP(3))) XOR ((OP(4) XOR OP(5)) XOR (OP(6) XOR OP(7))))
		XOR (((OP(8) XOR OP(9)) XOR (OP(10) XOR OP(11))) XOR ((OP(12) XOR OP(13)) XOR (OP(14) XOR OP(15))));
	SOM(1) <= (OP(1) XOR OP(3)) OR (OP(5) XOR OP(7)) OR (OP(9) XOR OP(11)) OR (OP(13) XOR OP(15));
		SOM(2) <= (OP(3) XOR OP(7)) OR (OP(11) XOR OP(15));
	SOM(3) <= OP(7) XOR OP(15);
	SOM(4) <= OP(15);

	Q_A(4) <= IN_KEYBOARD(16);

	ADD_SOM: SOMADOR8B PORT MAP(Q_A, SOM, '0', OUT_KEY, C_OUT);

END DECODING;